moudle test()    
    
    logic [3:0] D,
    logic clk, rst